library IEEE;
use IEEE.std_logic_1164.all;
use IEEE..all

entity 4to1Mux is 
  port( D0,D1,D2,D3:in std_logic;
       select: in std_logic 
